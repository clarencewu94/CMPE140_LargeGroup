module soc_addr_dec(
        input wire WE,
        input wire [31:0] A, // Check size
        output wire WE1,
        output wire WE2,
        output wire WEM,
        output wire [1:0] RdSel
    );

    


endmodule