module gpio(
        input wire clk,
        input wire reset,
        input wire [1:0] A,
        input wire WE2,
        input wire [31:0] WD,
        output wire RD
    );




endmodule